-- MCU Command Control (MCUCC) Component
-- Robotics Club at UCF
-- Jonathan Mohlenhoff - jmohlenh@ist.ucf.edu

library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;

use work.MCUPRT.all;
use work.mux2to1.all;
use work.rcOut.all;
use work.rcIn.all;
use work.ADC.all;
--use work.ADCSlow.all;
use work.SevenSegment.all;

entity mcuccComp is
	Port
	(
			TXD          : out std_logic;
			RXD          : in std_logic;
			clock        : in std_logic;
			d_out        : out std_logic_vector (7 downto 0) := x"00";
			d_in			 : in std_logic_vector (7 downto 0) := x"00";
			rc_out       : out std_logic_vector (7 downto 0); -- physical pins connected to motors
			rc_REMOTE : in std_logic_vector (7 downto 0);  --  signals passed to motors via mux
			
			--Pmod AD1 interface signals for battery
			ad0_SDATA0   : in std_logic;
			ad0_SDATA1   : in std_logic;
			ad0_SCLK     : out std_logic;
			ad0_nCS      : out std_logic;
			
			--Pmod AD1 interface signals for arm actuator
			ad1_SDATA0   : in std_logic;
			ad1_SDATA1   : in std_logic;
			ad1_SCLK     : out std_logic;
			ad1_nCS      : out std_logic;
			
			leds	       : out std_logic_vector (7 downto 0);
			switch		 : in std_logic_vector (7 downto 0);
			btn			 : in std_logic_vector (3 downto 0);
													
			sevenSegC	 : out std_logic_vector(6 downto 0);
			sevenSegA	 : out std_logic_vector(3 downto 0)
	);
end mcuccComp;

architecture Behavioral of mcuccComp is
	
	signal rt_commandRx : std_logic_vector (7 downto 0);
	signal rt_dataRx : std_logic_vector (31 downto 0);
	signal rt_packetRx : std_logic;
	signal rt_packetRd : std_logic;
	
	signal rt_commandTx : std_logic_vector (7 downto 0);
	signal rt_dataTx : std_logic_vector (31 downto 0);
	signal rt_packetTx : std_logic;
	signal rt_packetSent : std_logic; -- buffer is empty
	
	signal rc_outValue0 : std_logic_vector (7 downto 0) := x"80";  -- 
	signal rc_outValue1 : std_logic_vector (7 downto 0) := x"80";  --
	signal rc_outValue2 : std_logic_vector (7 downto 0) := x"80";  -- 
	signal rc_outValue3 : std_logic_vector (7 downto 0) := x"80";  --
	signal rc_outValue4 : std_logic_vector (7 downto 0) := x"80";  --
	signal rc_outValue5 : std_logic_vector (7 downto 0) := x"80";  --
	signal rc_outValue6 : std_logic_vector (7 downto 0) := x"80";  --
	signal rc_outValue7 : std_logic_vector (7 downto 0) := x"80";  --
	
	signal rc_outFPGA   : std_logic_vector (7 downto 0);  --  signals generated by FPGA as per computer's request
	
	signal rc_inValue0  : std_logic_vector (7 downto 0);  -- Value read from module to set signal mode
	signal rc_inValue1  : std_logic_vector (7 downto 0);  -- Value read from module to set signal mode
	signal rc_inValue2  : std_logic_vector (7 downto 0);  -- Value read from module to set signal mode
	signal rc_inValue3  : std_logic_vector (7 downto 0);  -- Value read from module to set signal mode
	signal rc_inValue4  : std_logic_vector (7 downto 0);  -- Value read from module to set signal mode
	signal rc_inValue5  : std_logic_vector (7 downto 0);  -- Value read from module to set signal mode
	signal rc_inValue6  : std_logic_vector (7 downto 0);  -- Value read from module to set signal mode	
	
	signal mode         : std_logic;                      -- signal to determine where boat control lies
																		   -- Computer, FPGA or Human
	signal rc_Count     : std_logic_vector (7 downto 0);
	
	type commandState is (waitForCommand, processCommand);
	signal commandStateCurrent : commandState := waitForCommand;
	signal commandStateNext : commandState;
	

	signal ad0_data0		: std_logic_vector (11 downto 0);
	signal ad0_data1		: std_logic_vector (11 downto 0);
	signal ad0_start		: std_logic;
	signal ad0_done		: std_logic;
	signal ad0_reset		: std_logic := '0';
	
	signal ad0_analog0	: std_logic_vector (11 downto 0);
	signal ad0_analog1	: std_logic_vector (11 downto 0);
	
	--Signals for linear actuator and pivot
	
	signal ad1_data0		: std_logic_vector (11 downto 0);
	signal ad1_data1		: std_logic_vector (11 downto 0);
	signal ad1_start		: std_logic;
	signal ad1_done		: std_logic;
	signal ad1_reset		: std_logic := '0';
	
	signal ad1_analog0	: std_logic_vector (11 downto 0);
	signal ad1_analog1	: std_logic_vector (11 downto 0);
	
	signal pivot_setpoint : std_logic_vector (7 downto 0) := x"80";
	signal linear_setpoint : std_logic_vector (7 downto 0) := x"00";
	
	signal digit0, digit1, digit2, digit3 : std_logic_vector(3 downto 0);

begin

	mcuprt_module: mcuprtComp port map
	(
		TXD => TXD,
		RXD => RXD,
		clock => clock,
		commandRx => rt_commandRx,
		dataRx => rt_dataRx,
		packetRx => rt_packetRx,
		packetRd => rt_packetRd,
		commandTx => rt_commandTx,
		dataTx => rt_dataTx,
		packetTx => rt_packetTx,
		packetSent => rt_packetSent
	);
	
	--Left Motor (Muxed by Transmitter Right Stick)
	rc_in0_module: rcInComp port map
	(
		rcIn => rc_REMOTE(0),
		rcValue => rc_inValue0,
		clock => clock
	);
	
	--Right Motor (Muxed by Transmitter Right Stick)
	rc_in1_module: rcInComp port map
	(
		rcIn => rc_REMOTE(1),
		rcValue => rc_inValue1,
		clock => clock
	);
	
	--Comp / RC Control (Left Stick Up/Down Value)
	rc_in2_module: rcInComp port map
	(
		rcIn => rc_REMOTE(2),
		rcValue => rc_inValue2,
		clock => clock
	);

	--Lateral (Left Stick Left/Right Value)
	rc_in3_module: rcInComp port map
	(
		rcIn => rc_REMOTE(3),
		rcValue => rc_inValue3,
		clock => clock
	);

	--ESTOP (Switch)
	rc_in4_module: rcInComp port map
	(
		rcIn => rc_REMOTE(4),
		rcValue => rc_inValue4,
		clock => clock
	);

	--Pump (Knob)
	rc_in5_module: rcInComp port map
	(
		rcIn => rc_REMOTE(5),
		rcValue => rc_inValue5,
		clock => clock
	);

	-- (Switch B)
	rc_in6_module: rcInComp port map
	(
		rcIn => rc_REMOTE(6),
		rcValue => rc_inValue6,
		clock => clock
	);
	
	rc_out0_module: rcOutComp port map
	(
		rcOut => rc_outFPGA(0),
		rcValue => rc_outValue0,
		clock => clock
	);
	 
	rc_out1_module: rcOutComp port map
	(
		rcOut => rc_outFPGA(1),
		rcValue => rc_outValue1,
		clock => clock
	);
	 
	rc_out2_module: rcOutComp port map
	(
		rcOut => rc_outFPGA(2),
		rcValue => rc_outValue2,
		clock => clock
	);
	 
	rc_out3_module: rcOutComp port map
  	(
		rcOut => rc_outFPGA(3),
		rcValue => rc_outValue3,
		clock => clock
	);
	 
	rc_out4_module: rcOutComp port map
	(
		rcOut => rc_outFPGA(4),
		rcValue => rc_outValue4,
		clock => clock
	 );
	 
	 rc_out5_module: rcOutComp port map
	(
		rcOut => rc_outFPGA(5),
		rcValue => rc_outValue5,
		clock => clock
	 );
	 
	 rc_out6_module: rcOutComp port map
	(
		rcOut => rc_outFPGA(6),
		rcValue => rc_outValue6,
		clock => clock
	 );
	 
	rc_out7_module: rcOutComp port map
	(
		rcOut => rc_outFPGA(7),
		rcValue => rc_outValue7,
		clock => clock
	 );
	 
	 --Left Motor
	 muxRC0_module: mux2to1Comp port map
	 (
		inputA => rc_outFPGA(0),
		inputB => rc_REMOTE(0),
		sel => mode,
		output => rc_out(0)
	 );
	 
	 --Right Motor
	 muxRC1_module: mux2to1Comp port map
	 (
		inputA => rc_outFPGA(1),
		inputB => rc_REMOTE(1),
		sel => mode,
		output => rc_out(1)
	 );
	 
	 --Lateral
	 muxRC2_module: mux2to1Comp port map
	 (
		inputA => rc_outFPGA(2), --Laterl channel from computer
		inputB => rc_REMOTE(3), --Lateral channel from transmitter
		sel => mode,
		output => rc_out(2) --Lateral channel to motor
	 );
	 
	 --Pump
	 muxRC3_module: mux2to1Comp port map
	 (
		inputA => rc_outFPGA(3),
		inputB => rc_REMOTE(5), --Knob on Transmitter
		sel => mode,
		output => rc_out(3)
	 );
	 
	 ad0: AD1RefComp port map
	 (
		  --General usage
		CLK => clock,      
		RST => ad0_reset, 
     
		--Pmod interface signals
		SDATA1 => ad0_SDATA0,
		SDATA2 => ad0_SDATA1,
		SCLK => ad0_SCLK,
		nCS => ad0_nCS,   
        
		--User interface signals
		 DATA1 => ad0_data0,
		 DATA2 => ad0_data1,
		 START => ad0_start,
		 DONE  => ad0_done
	 );
	 
	 ad1: AD1RefComp port map
	 (
		  --General usage
		CLK => clock,      
		RST => ad1_reset, 
     
		--Pmod interface signals
		SDATA1 => ad1_SDATA0,
		SDATA2 => ad1_SDATA1,
		SCLK => ad1_SCLK,
		nCS => ad1_nCS,   
        
		--User interface signals
		 DATA1 => ad1_data0,
		 DATA2 => ad1_data1,
		 START => ad1_start,
		 DONE  => ad1_done
	 );
	 
	 sevenSegment: SegmentRefComp port map
    (    
		CLK	 => clock,
		input1 => digit0,
		input2 => digit1,
		input3 => digit2,
		input4 => digit3,
		sevenseg1 => sevenSegC,
		anodes => sevenSegA
	);
	 
	 ad0_reset <= '0';
	 ad1_reset <= '0';
	 

	 --ALWAYS COMPUTER CONTROLLED
	 --pan
	 rc_out(4) <= rc_outFPGA(4);
	 
	 --Tilt
	 rc_out(5) <= rc_outFPGA(5);

	 --Arm_pivot
	 rc_out(6) <= rc_outFPGA(6);
	 
	 --Arm_linear
	 rc_out(7) <= rc_outFPGA(7);

	 --Comp / RC Control
	 --d_in(2) <= mode; 
	 d_out(7) <= mode;

	 --leds <= ad1_analog0 (11 downto 4);
	 
	 
process(clock)
	begin
		if (rising_edge(clock)) then
			commandStateCurrent <= commandStateNext;
		end if;
	end process;


--Controls Computer / RC Mode from Receiver's Channel 3 (Left Stick Up/Down)
process(clock)
	begin
		if(rising_edge(clock)) then
			if (rc_inValue2 < x"67") then
				mode <= '0';
			elsif (rc_inValue2 > x"98") then
				mode <= '1';
			else
				-- in hysterisis (do nothing)
			end if;
		end if;
end process;

process(clock, rt_commandRx)
	variable tempD_outPort, tempD_outValue: std_logic_vector (7 downto 0);
	variable servo_port   : std_logic_vector (7 downto 0);
	variable input_port : std_logic_vector (7 downto 0);
	variable input_value : std_logic_vector (7 downto 0);
	begin
		if (rising_edge(clock)) then
			if (commandStateCurrent = commandStateNext) then
				case commandStateCurrent is
					when waitForCommand =>
						rt_packetTx <= '0';
						if (rt_packetRx = '1') then
							rt_packetRd <= '1';
							commandStateNext <= processCommand;
						else
							commandStateNext <= waitForCommand;
						end if;
					
					when processCommand =>
						if (rt_packetSent = '1') then -- if a complete packet has been sent
							case rt_commandRx is
								when x"0D" => --Ping Message Received
									rt_commandTx <= x"84"; --Pong Command to be sent in respone
									rt_dataTx (7 downto 0) <= x"50";
									rt_dataTx (15 downto 8) <= x"4F";
									rt_dataTx (23 downto 16) <= x"4E";
									rt_dataTx  (31 downto 24) <= x"47";
									rt_packetTx <= '1'; -- ready to transmit
								
								when x"0C" => -- set Digital output message received
									tempD_outPort := rt_dataRx (7 downto 0);
									tempD_outValue := rt_dataRx (15 downto 8);
									case tempD_outPort is
										when x"00" =>
											d_out(0) <= tempD_outValue(0);
											
										when x"01" =>
											d_out(1) <= tempD_outValue(1);
										
										when x"02" =>  -- Outside BLUE LED for Comp/RC control
											d_out(2) <= tempD_outValue(2);
											
										when x"03" =>
											d_out(3) <= tempD_outValue(3);
										
										when x"04" =>
											d_out(4) <= tempD_outValue(4);
											
										when x"05" =>
											d_out(5) <= tempD_outValue(5);
											
										when x"06" =>
											d_out(6) <= tempD_outValue(6);
											
										--when x"07" =>
											--d_out(7) <= tempD_outValue(7);	
										
										when others =>
											-- port not defined
									end case;
								
								when x"0B" => -- Set Servo Out Message Received
									servo_port := rt_dataRx (7 downto 0);
									--sValue_out <= rt_dataRx (15 downto 8);
									
									case servo_port is 
										when x"00" => -- Left Motor
											rc_outValue0 <= rt_dataRx (15 downto 8);
											
										when x"01" => -- Right Motor
											rc_outValue1 <= rt_dataRx (15 downto 8);
											
										when x"02" => -- Lateral Motor
											rc_outValue2 <= rt_dataRx (15 downto 8);
											
										when x"03" => -- Pump
											rc_outValue3 <= rt_dataRx (15 downto 8);
											
										when x"04" => -- Pan
											rc_outValue4 <= rt_dataRx (15 downto 8);
										
										when x"05" => -- Tilt
											rc_outValue5 <= rt_dataRx (15 downto 8);
											
										when x"06" => -- Arm Pivot
											pivot_setpoint <= rt_dataRx (15 downto 8);
											--rc_outValue6 <= rt_dataRx (15 downto 8);
											
										when x"07" => -- Arm Linear
											--linear_setpoint <= rt_dataRx (15 downto 8);
											rc_outValue7 <= rt_dataRx (15 downto 8);
										when others =>
											-- do nothing fool
									end case;
								
								when x"82" => --Report Digital Input Message Received
									case rt_dataRx (7 downto 0) is
										when x"00" => -- Port 0 Inputs
											input_value := d_in;

										when others =>
											--Invalid port received
											input_value := x"00";
									end case;
									
									rt_commandTx <= x"82"; --Report Digital Input
									rt_dataTx (7 downto 0) <= rt_dataRx (7 downto 0);
									rt_dataTx (15 downto 8) <= input_value;
									rt_dataTx (23 downto 16) <= x"00";
									rt_dataTx  (31 downto 24) <= x"00";
									rt_packetTx <= '1'; -- ready to transmit
									
								when x"83" =>
									case rt_dataRx (7 downto 0) is
										when x"00" =>
											rt_commandTx <= x"83"; --Report Analog Input
											rt_dataTx (7 downto 0) <= x"00";
											rt_dataTx (23 downto 8) <= x"0" & ad0_analog0; --Batt Motors
											rt_dataTx  (31 downto 24) <= x"00";
											rt_packetTx <= '1'; -- ready to transmit
										
										when x"01" =>
											rt_commandTx <= x"83"; --Report Analog Input
											rt_dataTx (7 downto 0) <= x"01";
											rt_dataTx (23 downto 8) <= x"0" & ad0_analog1; --Batt Electronics
											rt_dataTx  (31 downto 24) <= x"00";
											rt_packetTx <= '1'; -- ready to transmit
											
										when x"02" =>
											rt_commandTx <= x"83"; --Report Analog Input
											rt_dataTx (7 downto 0) <= x"02";
											rt_dataTx (23 downto 8) <= x"0" & ad1_analog0; --Pivot Arm
											rt_dataTx  (31 downto 24) <= x"00";
											rt_packetTx <= '1'; -- ready to transmit
										
										when x"03" =>
											rt_commandTx <= x"83"; --Report Analog Input
											rt_dataTx (7 downto 0) <= x"03";
											rt_dataTx (23 downto 8) <= x"0" & ad1_analog1; --Arm Extension
											rt_dataTx  (31 downto 24) <= x"00";
											rt_packetTx <= '1'; -- ready to transmit
										
										when others =>
											--Invalid analog port
									end case;
								
								when x"88" => --Report Servo Input Message Received
									case rt_dataRx (7 downto 0) is
										when x"00" => -- start button status
											rt_dataTx (15 downto 8) <= rc_inValue0;
											
										when x"01" =>
											rt_dataTx (15 downto 8) <= rc_inValue1;
										
										when x"02" =>
											rt_dataTx (15 downto 8) <= rc_inValue2;
										
										when x"03" =>
											rt_dataTx (15 downto 8) <= rc_inValue3;
										
										when x"04" =>
											rt_dataTx (15 downto 8) <= rc_inValue4;
										
										when x"05" =>
											rt_dataTx (15 downto 8) <= rc_inValue5;
										
										when x"06" =>
											rt_dataTx (15 downto 8) <= rc_inValue6;
										
										when others =>
											--Invalid channel received
									end case;									
								
									rt_commandTx <= x"88"; --Report Servo Input
									rt_dataTx (7 downto 0) <= rt_dataRx (7 downto 0);
									rt_dataTx (23 downto 16) <= x"00";
									rt_dataTx  (31 downto 24) <= x"00";
									rt_packetTx <= '1'; -- ready to transmit
								
								when others =>
									
							end case;
							commandStateNext <= waitForCommand;
							
						else
							rt_packetTx <= '0';
						end if;
					
				end case;
			end if;
		end if;
	end process;
	
ad0_process: process(clock)
	
	begin
	
		if (rising_edge(clock)) then
			if (ad0_done = '1') then
				ad0_analog0 <= ad0_data0;
				ad0_analog1 <= ad0_data1;
				ad0_start <= '1';
			else
				ad0_start <= '0';
			end if;
		end if;
	
	end process;
	
ad1_process: process(clock)
	type table is array (0 to 127) of std_logic_vector (23 downto 0);
	variable movingAverageTable1 : table;
	variable movingAverageTable2 : table;
	variable doneCount : integer := 0;
	variable tempAverage1 : std_logic_vector (23 downto 0) := x"000000";
	variable tempAverage2 : std_logic_vector (23 downto 0) := x"000000";
	
	begin
	
		if (rising_edge(clock)) then
			if (ad1_done = '1') then
				ad1_analog0 <= ad1_data0;
				ad1_analog1 <= ad1_data1;
				
--				tempAverage1 := tempAverage1 - movingAverageTable1(doneCount);
--				tempAverage2 := tempAverage2 - movingAverageTable2(doneCount);
--				movingAverageTable1(doneCount) := x"000" & ad1_data0;
--				movingAverageTable2(doneCount) := x"000" & ad1_data1;
--				tempAverage1 := tempAverage1 + movingAverageTable1(doneCount);
--				tempAverage2 := tempAverage2 + movingAverageTable2(doneCount);
--				
--				doneCount := doneCount + 1;
--				if (doneCount > 15) then
--					doneCount := 0;
--				end if;
--				
--				ad1_analog0 <= tempAverage1 (18 downto 7);
--				ad1_analog1 <= tempAverage2 (18 downto 7);
				
				ad1_start <= '1';
			else
				ad1_start <= '0';
			end if;
		end if;
	
	end process;

--
--linear_control: process(clock)
--variable linear_position: std_logic_vector (7 downto 0);
--variable hyst_state: std_logic := '0';
--variable small_window : std_logic_vector (7 downto 0) := x"08";
--variable big_window : std_logic_vector (7 downto 0) := x"20";
--variable linear_setpoint_temp : std_logic_vector (7 downto 0);
--variable hyst_counter_high : integer := 0;
--variable hyst_counter_low : integer := 0;
--variable hyst_counter_limit : integer := 2048;
--	begin
--		if (rising_edge(clock) and (ad1_done = '1')) then
--			linear_position := ad1_analog1 (11 downto 4);
--			
--			if (hyst_state = '0') then
--				if (linear_setpoint < small_window) then
--					linear_setpoint_temp := small_window;
--				elsif (linear_setpoint > (x"FF" - small_window)) then
--					linear_setpoint_temp := x"FF" - small_window;
--				else
--					linear_setpoint_temp := linear_setpoint;
--				end if;
--				
--				if (linear_position < linear_setpoint_temp - small_window) then 
--					hyst_counter_low := 0;
--					hyst_counter_high := 0;
--					--rc_outValue7 <= x"FF";
--					
--				elsif (linear_position > linear_setpoint_temp + small_window) then
--					hyst_counter_low := 0;
--					hyst_counter_high := 0;
--					--rc_outValue7 <= x"00";
--					
--				else
--					--rc_outValue7 <= x"80";
--					hyst_counter_high :=	hyst_counter_high + 1;
--					if (hyst_counter_high > hyst_counter_limit) then
--						hyst_counter_high := 0;
--						hyst_counter_low := 0;
--						hyst_state := '1';
--					end if;
--				end if;
--	
--			else
--				if (linear_setpoint < big_window) then
--					linear_setpoint_temp := big_window;
--				elsif (linear_setpoint > (x"FF" - big_window)) then
--					linear_setpoint_temp := x"FF" - big_window;
--				else
--					linear_setpoint_temp := linear_setpoint;
--				end if;
--				
--    			if (linear_position < (linear_setpoint_temp - big_window)) then 
--					hyst_counter_high := 0;
--					hyst_counter_low := hyst_counter_low + 1;
--					if (hyst_counter_low > hyst_counter_limit) then
--						hyst_counter_low := 0;
--						hyst_counter_high := 0;
--						hyst_state := '0';
--					end if;
--					
--				elsif (linear_position > (linear_setpoint_temp + big_window)) then
--					hyst_counter_low := 0;
--					hyst_counter_high := hyst_counter_high + 1;
--					if (hyst_counter_high > hyst_counter_limit) then
--						hyst_counter_low := 0;
--						hyst_counter_high := 0;
--						hyst_state := '0';
--					end if;
--					
--				else
--					--rc_outValue7 <= x"80";
--					hyst_counter_high := 0;
--					hyst_counter_low := 0;
--				end if;
--			
--			end if;
--			
--		end if;
--	end process;
	
pivot_pid: process(clock)
	variable p : signed(31 downto 0) := to_signed(3, 32);
	variable i : signed(31 downto 0) := to_signed(0, 32);
	variable d : signed(31 downto 0) := to_signed(15, 32);
	variable desiredSetpoint : signed(31 downto 0) := to_signed(0, 32);
	variable currentSetpoint : signed(31 downto 0) := to_signed(0, 32);
	variable position : signed(31 downto 0) := to_signed(0, 32);
	variable error : signed(31 downto 0) := to_signed(0, 32);
	variable previousError : signed(31 downto 0) := to_signed(0, 32);
	variable errorSum : signed(31 downto 0) := to_signed(0, 32);
	variable output : signed(31 downto 0) := to_signed(0, 32);
	variable offset : signed(31 downto 0) := to_signed(128, 32);
	variable counter : signed(31 downto 0) := to_signed(0, 32);
	variable period : signed(31 downto 0) := to_signed(1000000, 32);
	variable display : std_logic_vector(31 downto 0);
	variable absErrorSum : signed(31 downto 0) := to_signed(0, 32);
	begin
		if(rising_edge(clock)) then
			counter := counter + to_signed(1, 32);
			if(counter > period) then
				counter := to_signed(0, 32);
				
				--p := signed(x"0000000" & switch (3 downto 0));
				--i := signed(x"0000000" & switch (7 downto 4));
				--d := signed(x"0000000" & switch (7 downto 4));
				
				
				--position := x"00000080";
				--setpoint := x"0000007F";
				position := signed(x"000000" & ad1_analog0 (11 downto 4));
				desiredSetpoint := signed(x"000000" & pivot_setpoint);
				
				--Ramp the desired setpoint
				if (desiredSetpoint > currentSetpoint) then
					currentSetpoint := currentSetpoint + to_signed(1, 32);
					if (currentSetpoint > desiredSetpoint) then
						currentSetpoint := desiredSetpoint;
					end if;
				
				elsif (desiredSetpoint < currentSetpoint) then
					currentSetpoint := currentSetpoint - to_signed(1, 32);
					if (currentSetpoint < desiredSetpoint) then
						currentSetpoint := desiredSetpoint;
					end if;
				end if;
				
				previousError := error;
				error := currentSetpoint - position;
				output := p*error + i*errorSum/2 + d*(error - previousError) + offset;
			
				if (output < to_signed(0, 32)) then
					output := to_signed(0, 32);
				elsif (output > to_signed(255, 32)) then
					output := to_signed(255, 32);
				else
					--errorSum := errorSum + error;
				end if;
				
--				if (btn(1 downto 0) = "00") then
--					if (errorSum < to_signed(0, 32)) then
--						leds(0) <= '1';
--					else
--						leds(0) <= '0';
--					end if;
--					absErrorSum := abs(errorSum);
--					display := std_logic_vector(absErrorSum);
--				elsif (btn(1 downto 0) = "01") then
--					if (error < to_signed(0, 32)) then
--						leds(0) <= '1';
--					else
--						leds(0) <= '0';
--					end if;
--					absErrorSum := abs(error);
--					display := std_logic_vector(absErrorSum);
--				elsif (btn(1 downto 0) = "10") then
--					if (output < to_signed(0, 32)) then
--						leds(0) <= '1';
--					else
--						leds(0) <= '0';
--					end if;
--					absErrorSum := abs(output);
--					display := std_logic_vector(absErrorSum);
--				end if;
--				
--				digit0 <= display (3 downto 0);
--				digit1 <= display (7 downto 4);
--				digit2 <= display (11 downto 8);
--				digit3 <= display (15 downto 12);
				
				rc_outValue6 <= std_logic_vector(output(7 downto 0));				
			end if;
		end if;
	end process;

end Behavioral;

